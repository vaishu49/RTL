// Code your design here

module not_dut(y,a);
  input a;
  output y;
  assign  y = ~a;
  
endmodule
